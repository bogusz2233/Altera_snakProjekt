
module unsaved (
	clkout_clk,
	clk_in_clk,
	reset_reset);	

	output		clkout_clk;
	input		clk_in_clk;
	input		reset_reset;
endmodule
