LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;


ENTITY READING IS 
PORT(
		CLK 		:IN 	STD_LOGIC;							-- CLK = 100 ms;
		ODCZYT	:OUT 	STD_LOGIC_VECTOR(7 DOWNTO 0); -- DO CENTRAL UNIT
		
		CMD		:OUT 	STD_LOGIC_VECTOR(7 DOWNTO 0);	--	ROZKAZ DLA SHIFT
		CLKSHIFT :OUT	STD_LOGIC;							-- DO TAKTOWANIA SHIFTA
		DATA		:IN 	STD_LOGIC_VECTOR(7 DOWNTO 0);	--ODCZYT ZE SFITHA
		TRANS		:IN	STD_LOGIC;
);
END READING;

ARCHITECTURE MAIN OF READING IS 
	/*
	SETUP - POCZATEK USTAWIENIE POCZATKOWE , POWROT DO TEGO STANU PO KAŻDY SKONCZONYM ODZCZYCIE
	ASK	- WYSLANIE PRZEZ SHIFT INFORMACJI ZE PROSI O  KOMUNIKACJE
	BEGINCOM		-	WYSLANIE PRZEZ SHIFT INFORMACJI ŻE  PROSI O ODCZYT
	FIRSTREAD	-	PIERWSZY ODCZYT (NIC TUTAJ NIE CZYTA)
	DIRREAD		- CZYTA TUTAJ STRZALKI KONTROLERA 
	*/
	TYPE STANY 				IS (SETUP,ASK,BEGINCOM,FIRREAD,DIRREAD) :=SETUP;
	SIGNAL ZEGAR : STD_LOGIC:=0;
	BEGIN
	
	CLKSHIFT<=ZEGAR;
	
	PROCESS(CLK)
		BEGIN 
		IF RISING_EDGE (CLK)
			ZEGAR<= NOT ZEGAR;
			CASE STANY IS
				WHEN SETUP =>
					CMD=OTHERS(=>'0');
					ODCZYT <=DATA;
				WHEN ASK =>
					IF TRANS='1' THEN
						CMD<="0000_0001";
					ELSE 
						STAN :=BEGINCOM;
					END IF;
				WHEN BEGINCOM =>
					IF TRANS='1' THEN
						CMD<="0100_0010";
					ELSE 
						STAN :=FIRREAD;
					END IF;
				WHEN FIRREAD=>
					IF TRANS='1' THEN
						CMD<="1111_1111";
					ELSE 
						STAN :=DIRREAD;
					END IF;
				WHEN DIRREAD=>
					IF TRANS='1' THEN
						CMD<="1111_1111";
					ELSE 
						STAN :=SETUP;
					END IF;
				
			END CASE;
		END IF;
	END PROCESS;
END MAIN;