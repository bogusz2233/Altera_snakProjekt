LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

ENTITY SHIFT IS 
	PORT(
			CLK 		: IN STD_LOGIC; 							--ZEGAR Z READ
			CMD_IN 	: IN STD_LOGIC_VECTOR(7 DOWNTO 0);	--KOMENDA Z READ
			DATA		: IN STD_LOGIC;							-- ZCZYTANIE WARTOSCI Z PINU
			ODCZYT	: OUT STD_LOGIC_VECTOR(7 DOWTO 0);
			CMDPIN	: OUT STD_LOGIC;
			TRANS		: OUT STD_LOGIC;	-- DO STEROWANIA READ'EM
	);

END SHIFT;

ARCHITECTURE MAIN OF SHIFT IS 

	TYPE STANY IS (WAITING,SENDCMD,READDA, PRINT):= WAITING
	SIGNAL LICZNIKBIT	:INTEGER RANGE 0 TO 8:=0;
	SIGNAL ZCZYTANIE	:STD_LOGIC_VECTOR(7 DOWTO 0);

	BEGIN
	PROCESS(CLK)
		IF RISING_EDGE (CLK)
			CASE STANY IS
				WHEN WAITING =>
					IF(CMD_IN)<="0000_0000") THEN
						STANY :=WAITING;
					ELSE
						STANY := SENDCMD
						LICZNIKBIT:=0;
						TRANS <='1';
					END IF;
				WHEN SENDCMD=>
					IF LICZNIKBIT >7 THEN 
						LICZNIKBIT = 0;
						STANY :=READDA;
					END IF;
					CMDPIN<=CMD_IN(LICZNIKBIT );
					LICZNIKBIT := LICZNIKBIT + 1;
				WHEN READDA =>
					IF LICZNIKBIT >7 THEN 
						LICZNIKBIT = 0;
						STANY := PRINT;
					END IF;
					ZCZYTANIE(LICZNIKBIT ) <= DATA;
					LICZNIKBIT := LICZNIKBIT + 1;
				WHEN PRINT =>
					ODCZYT <= ZCZYTANIE;
					TRANS <='0';
					STANY :=WAITING;
		END IF;
	END PROCESS;
END MAIN;