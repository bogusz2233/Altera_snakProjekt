LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

ENTITY Controller_PS1 IS 
PORT(
		-- PIN CONNECTED TO CONTROLLER	  \/ TO CONNECT
		DATA_PIN		:IN STD_LOGIC;			-- 1 PIN		-- PULL_UP;
		CMD_PIN		:OUT STD_LOGIC;		--	2 PIN
		ATT_PIN		:OUT STD_LOGIC;		--	6 PIN
		CLOCK_PIN	:OUT STD_LOGIC;		--	7 PIN	 	-- REATING AT FALLING EDGE
											--GND -- 4 PIN
									--VCC(3,3V)	--	5 PIN
		CLK			:IN STD_LOGIC;							-- REATING AT RISING_EDGE
);	
END Controller_PS1;

ARCHITECTURE MAIN OF Controller_PS1 IS

	TYPE STANY 				IS (SETUP,READING) :=SETUP;
	
	SIGNAL DATA,CMD, ATT,CLOCK;
	BEGIN
	-- ASSIGNING INSIDE STATE  TO PIN
	CMD_PIN <= CMD;
	ATT_PIN <= ATT;
	CLOCK_PIN <= CLOCK;
	
	PROCESS(CLK)
		BEGIN 
		IF RISING_EDGE (CLK)
		CASE STANY IS
			WHEN SETUP =>
				ATT <= '1';
				CLOCK <= '1';
			WHEN READING =>
				ATT<='0'
				
			
	END PROCESS;
END MAIN;