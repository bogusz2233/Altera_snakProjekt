LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

ENTITY SYNC_640x480 IS
PORT(
	CLK_25MHz		: IN STD_LOGIC;
	-- DO SYNCHRONIZACJI I DO WYSTAWIENIA CZARNEGO KOLORU GDY SĄ PUSTE  PIKSELE
	HSYNC,VSYNC 	: OUT STD_LOGIC;
	BLACK				: OUT STD_LOGIC;
	
	-- DO CENTRALI, DZIEKI TEMU BĘDZIE MOGŁA SIE ONA SYNCHRONIZOWAĆ Z WYSWIETLACZEM
	HPOS_OUT			: OUT STD_LOGIC_VECTOR(10 DOWNTO 0);
	VPOS_OUT			: OUT STD_LOGIC_VECTOR(10 DOWNTO 0)
);


END ENTITY;

ARCHITECTURE MAIN OF SYNC_640x480 IS
	
	-- OBECNY PIKSEL
	SIGNAL HPOS			:INTEGER RANGE 0 TO 800	:=0; 
	SIGNAL VPOS			:INTEGER RANGE 0 TO 524	:=0;
	SIGNAL EMPTY 		:STD_LOGIC;		-- DO OKREŚLANIA CZY TERAZ SĄ PUSTE KOLORY 

		
	
	BEGIN
	BLACK <= EMPTY;

	PROCESS(CLK_25MHz)
	
	BEGIN
		
		IF(CLK_25MHz'EVENT AND CLK_25MHz ='1') THEN
			--PRZESŁANIE WIADOŚCI O POŁOŻENIU DO CENTRALNEGO UKŁADU
			IF(EMPTY = '0') THEN
				VPOS_OUT <= STD_LOGIC_VECTOR(TO_UNSIGNED(VPOS - 44 , VPOS_OUT'LENGTH) );
				HPOS_OUT	<= STD_LOGIC_VECTOR(TO_UNSIGNED(HPOS - 160, HPOS_OUT'LENGTH) ); 
				-- ODEJMUJE PUSTE BITY ŻEBY MIEĆ BEZWGLĘDNE POŁOŻENIA OBIEKTÓW
			END IF;

			IF(HPOS < 800) THEN
				HPOS<=HPOS + 1;
				ELSE
					--ZAKONCZENIE LINII
					HPOS<=0;
					IF(VPOS<524) THEN
					-- PRZESKOCZENIE DO NASTEPNIEJ LINNI
					VPOS<= VPOS + 1;
					ELSE
					-- ZAKONCZENIE RAMKI
					VPOS<=0;
				END IF;
			END IF;
			
			
			IF(HPOS > 16 AND HPOS< 112) THEN
				HSYNC<= '0';
				--EMPTY FRAME
			ELSE
				HSYNC<=	'1';
			END IF;
			
			IF(VPOS > 0 AND VPOS <13) THEN
				VSYNC <='0';
			ELSE 
				VSYNC <='1';
			END IF;
			
			IF((HPOS >0 AND HPOS< 160) OR (VPOS>0 AND VPOS <44)) THEN
					EMPTY <='1';
			ELSE 
					EMPTY <='0';
			END IF;
			
		END IF;
		END PROCESS;
		
	END ARCHITECTURE;
			