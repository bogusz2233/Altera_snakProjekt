LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY PLAYER_CONTROLER IS
PORT(
		UP_IN,DOWN_IN,LEFT_IN,RIGHT_IN 	: IN STD_LOGIC;
		UP,DOWN,LFT,RGT						: OUT STD_LOGIC;
		CLK_50HZ									: IN STD_LOGIC
);

END PLAYER_CONTROLER;

ARCHITECTURE MAIN OF PLAYER_CONTROLER IS
	BEGIN
		UP<= NOT UP_IN;
		DOWN<= NOT DOWN_IN;
		LFT<= NOT LEFT_IN;
		RGT<= NOT RIGHT_IN;
END MAIN;