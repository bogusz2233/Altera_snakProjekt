library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


PACKAGE FUNCTIONS IS
FUNCTION WYS_TO_LOGIC (ALL_P,PLACE_B, PLACE_E,POSITION, RESOLUTION :INTEGER) return INTEGER; --THIS FUNCTION CONVERT TO LOGIC POSION 

END PACKAGE;

PACKAGE BODY FUNCTIONS IS 

FUNCTION WYS_TO_LOGIC (ALL_P,PLACE_B, PLACE_E,POSITION,RESOLUTION :INTEGER) return INTEGER IS
	BEGIN
	RETURN (ALL_P -(POSITION -(PLACE_E - PLACE_B)) ) / RESOLUTION; 
	
END WYS_TO_LOGIC;
	
END PACKAGE BODY;