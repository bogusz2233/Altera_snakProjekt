LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY COLOR_STER IS 
PORT(
	BLACK_IN				: IN STD_LOGIC;
	RGB_IN				: IN STD_LOGIC_VECTOR(2 DOWNTO 0);
	R,G,B					: OUT STD_LOGIC
	);
END ENTITY;

ARCHITECTURE MAIN OF COLOR_STER IS

	BEGIN
	WITH BLACK_IN SELECT
	R <= RGB_IN(2) WHEN '0',
				'0' WHEN '1';
				
	WITH BLACK_IN SELECT
	G <= RGB_IN(1) WHEN '0',
				'0' WHEN '1';
	WITH BLACK_IN SELECT
	B <= RGB_IN(0) WHEN '0',
				'0' WHEN '1';
	

END MAIN;