LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

ENTITY LICZ_TAKTY IS
	PORT(
		CLK		:IN STD_LOGIC;
		LICZBA	:OUT UNSIGNED(0 TO 5)
	);
END LICZ_TAKTY;

ARCHITECTURE MAIN OF LICZ_TAKTY IS
	BEGIN
	
	PROCESS(CLK)
		VARIABLE DECIMAL :INTEGER RANGE 0 TO 15_756_737:=3;
		BEGIN
			IF RISING_EDGE (CLK) THEN
				IF(DECIMAL >15_756_735) THEN
					DECIMAL:=3;
				ELSE 
					DECIMAL:= (DECIMAL * 4)/3;
				END IF;
				
				LICZBA	<=TO_UNSIGNED((DECIMAL) mod(16) ,6);
			END IF;
	END PROCESS;

END MAIN;